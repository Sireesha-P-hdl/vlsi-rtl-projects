// Alarm Clock RTL Design
module alarm_clock();
endmodule
